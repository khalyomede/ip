
module ip

pub struct Ipv4 {
    pub mut:
        address [4]u8
}
