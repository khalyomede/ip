module ip

pub struct Ipv6 {
    pub mut:
        address [8]u16
}
