module ip

pub type Address = Ipv4 | Ipv6
